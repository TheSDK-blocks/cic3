../../../TheSDK_generators/verilog/cic3.v