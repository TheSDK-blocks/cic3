../../../TheSDK_generators/verilog/tb_cic3.v